module Hello(
    input a,
    output b
);
    assign b = a;
endmodule